// testcore.v

// Generated using ACDS version 14.0 209 at 2014.11.16.01:22:33

`timescale 1 ps / 1 ps
module testcore (
		input  wire        clk100_clk,            //         clk100.clk
		input  wire        reset_reset_n,         //          reset.reset_n
		output wire        led_export,            //            led.export
		input  wire        clk40_clk,             //          clk40.clk
		output wire [12:0] sdr_addr,              //            sdr.addr
		output wire [1:0]  sdr_ba,                //               .ba
		output wire        sdr_cas_n,             //               .cas_n
		output wire        sdr_cke,               //               .cke
		output wire        sdr_cs_n,              //               .cs_n
		inout  wire [15:0] sdr_dq,                //               .dq
		output wire [1:0]  sdr_dqm,               //               .dqm
		output wire        sdr_ras_n,             //               .ras_n
		output wire        sdr_we_n,              //               .we_n
		input  wire        adc_pll_locked_export, // adc_pll_locked.export
		output wire        mmc_nCS,               //            mmc.nCS
		output wire        mmc_SCK,               //               .SCK
		output wire        mmc_SDO,               //               .SDO
		input  wire        mmc_SDI,               //               .SDI
		input  wire        mmc_CD,                //               .CD
		input  wire        mmc_WP,                //               .WP
		input  wire        vga_clk,               //            vga.clk
		output wire [4:0]  vga_rout,              //               .rout
		output wire [4:0]  vga_gout,              //               .gout
		output wire [4:0]  vga_bout,              //               .bout
		output wire        vga_hsync_n,           //               .hsync_n
		output wire        vga_vsync_n,           //               .vsync_n
		output wire        vga_enable             //               .enable
	);

	wire         nios2_gen2_f_custom_instruction_master_multi_readra;                             // nios2_gen2_f:A_ci_multi_readra -> nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_readra
	wire         nios2_gen2_f_custom_instruction_master_multi_readrb;                             // nios2_gen2_f:A_ci_multi_readrb -> nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_readrb
	wire   [7:0] nios2_gen2_f_custom_instruction_master_multi_n;                                  // nios2_gen2_f:A_ci_multi_n -> nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_n
	wire         nios2_gen2_f_custom_instruction_master_done;                                     // nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_done -> nios2_gen2_f:A_ci_multi_done
	wire         nios2_gen2_f_custom_instruction_master_clk_en;                                   // nios2_gen2_f:A_ci_multi_clk_en -> nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_clken
	wire         nios2_gen2_f_custom_instruction_master_multi_writerc;                            // nios2_gen2_f:A_ci_multi_writerc -> nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_writerc
	wire  [31:0] nios2_gen2_f_custom_instruction_master_multi_result;                             // nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_result -> nios2_gen2_f:A_ci_multi_result
	wire         nios2_gen2_f_custom_instruction_master_clk;                                      // nios2_gen2_f:A_ci_multi_clock -> nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_clk
	wire         nios2_gen2_f_custom_instruction_master_reset_req;                                // nios2_gen2_f:A_ci_multi_reset_req -> nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire   [4:0] nios2_gen2_f_custom_instruction_master_multi_c;                                  // nios2_gen2_f:A_ci_multi_c -> nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_c
	wire   [4:0] nios2_gen2_f_custom_instruction_master_multi_b;                                  // nios2_gen2_f:A_ci_multi_b -> nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] nios2_gen2_f_custom_instruction_master_multi_a;                                  // nios2_gen2_f:A_ci_multi_a -> nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_a
	wire  [31:0] nios2_gen2_f_custom_instruction_master_multi_dataa;                              // nios2_gen2_f:A_ci_multi_dataa -> nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         nios2_gen2_f_custom_instruction_master_start;                                    // nios2_gen2_f:A_ci_multi_start -> nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_start
	wire  [31:0] nios2_gen2_f_custom_instruction_master_multi_datab;                              // nios2_gen2_f:A_ci_multi_datab -> nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_datab
	wire         nios2_gen2_f_custom_instruction_master_reset;                                    // nios2_gen2_f:A_ci_multi_reset -> nios2_gen2_f_custom_instruction_master_translator:ci_slave_multi_reset
	wire  [31:0] nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_result;        // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_result
	wire   [4:0] nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_b;             // nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_b -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_b
	wire   [4:0] nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_c;             // nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_c -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_c
	wire   [4:0] nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_a;             // nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_a -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_a
	wire         nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_clk_en;        // nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_clken -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire         nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_done;          // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_n;             // nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_n -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_n
	wire         nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_writerc;       // nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_clk;           // nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_clk -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_reset_req;     // nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_reset_req -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_start;         // nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_start -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_start
	wire  [31:0] nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_dataa;         // nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_readra;        // nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_readra -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire         nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_reset;         // nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_reset -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire  [31:0] nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_datab;         // nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_datab -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire         nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_readrb;        // nios2_gen2_f_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire  [31:0] nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_result;         // nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_result
	wire   [4:0] nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_b;              // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire   [4:0] nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_c;              // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_done;           // nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_done
	wire         nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire   [4:0] nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_a;              // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [7:0] nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_n;              // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire         nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_clk;            // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire         nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_start;          // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire  [31:0] nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_readra;         // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire         nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_reset;          // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire  [31:0] nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_datab;          // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire         nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire         nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // nios2_gen2_f_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire  [31:0] nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_result; // pixelsimd:result -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_start;  // nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_master_start -> pixelsimd:start
	wire  [31:0] nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> pixelsimd:dataa
	wire         nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_done;   // pixelsimd:done -> nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire         nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_master_clken -> pixelsimd:clk_en
	wire   [2:0] nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_n;      // nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_master_n -> pixelsimd:n
	wire         nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_master_reset -> pixelsimd:reset
	wire  [31:0] nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_master_datab -> pixelsimd:datab
	wire         nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // nios2_gen2_f_custom_instruction_master_multi_slave_translator0:ci_master_clk -> pixelsimd:clk
	wire         nios2_gen2_f_instruction_master_waitrequest;                                     // mm_interconnect_0:nios2_gen2_f_instruction_master_waitrequest -> nios2_gen2_f:i_waitrequest
	wire  [27:0] nios2_gen2_f_instruction_master_address;                                         // nios2_gen2_f:i_address -> mm_interconnect_0:nios2_gen2_f_instruction_master_address
	wire         nios2_gen2_f_instruction_master_read;                                            // nios2_gen2_f:i_read -> mm_interconnect_0:nios2_gen2_f_instruction_master_read
	wire  [31:0] nios2_gen2_f_instruction_master_readdata;                                        // mm_interconnect_0:nios2_gen2_f_instruction_master_readdata -> nios2_gen2_f:i_readdata
	wire         nios2_gen2_f_instruction_master_readdatavalid;                                   // mm_interconnect_0:nios2_gen2_f_instruction_master_readdatavalid -> nios2_gen2_f:i_readdatavalid
	wire         nios2_gen2_f_data_master_waitrequest;                                            // mm_interconnect_0:nios2_gen2_f_data_master_waitrequest -> nios2_gen2_f:d_waitrequest
	wire  [31:0] nios2_gen2_f_data_master_writedata;                                              // nios2_gen2_f:d_writedata -> mm_interconnect_0:nios2_gen2_f_data_master_writedata
	wire  [28:0] nios2_gen2_f_data_master_address;                                                // nios2_gen2_f:d_address -> mm_interconnect_0:nios2_gen2_f_data_master_address
	wire         nios2_gen2_f_data_master_write;                                                  // nios2_gen2_f:d_write -> mm_interconnect_0:nios2_gen2_f_data_master_write
	wire         nios2_gen2_f_data_master_read;                                                   // nios2_gen2_f:d_read -> mm_interconnect_0:nios2_gen2_f_data_master_read
	wire  [31:0] nios2_gen2_f_data_master_readdata;                                               // mm_interconnect_0:nios2_gen2_f_data_master_readdata -> nios2_gen2_f:d_readdata
	wire         nios2_gen2_f_data_master_debugaccess;                                            // nios2_gen2_f:jtag_debug_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_f_data_master_debugaccess
	wire         nios2_gen2_f_data_master_readdatavalid;                                          // mm_interconnect_0:nios2_gen2_f_data_master_readdatavalid -> nios2_gen2_f:d_readdatavalid
	wire   [3:0] nios2_gen2_f_data_master_byteenable;                                             // nios2_gen2_f:d_byteenable -> mm_interconnect_0:nios2_gen2_f_data_master_byteenable
	wire   [9:0] vga_m1_burstcount;                                                               // vga:avm_m1_burstcount -> mm_interconnect_0:vga_m1_burstcount
	wire         vga_m1_waitrequest;                                                              // mm_interconnect_0:vga_m1_waitrequest -> vga:avm_m1_waitrequest
	wire  [31:0] vga_m1_address;                                                                  // vga:avm_m1_address -> mm_interconnect_0:vga_m1_address
	wire         vga_m1_read;                                                                     // vga:avm_m1_read -> mm_interconnect_0:vga_m1_read
	wire  [31:0] vga_m1_readdata;                                                                 // mm_interconnect_0:vga_m1_readdata -> vga:avm_m1_readdata
	wire         vga_m1_readdatavalid;                                                            // mm_interconnect_0:vga_m1_readdatavalid -> vga:avm_m1_readdatavalid
	wire         mm_interconnect_0_nios2_gen2_f_debug_mem_slave_waitrequest;                      // nios2_gen2_f:jtag_debug_slave_waitrequest -> mm_interconnect_0:nios2_gen2_f_debug_mem_slave_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_gen2_f_debug_mem_slave_writedata;                        // mm_interconnect_0:nios2_gen2_f_debug_mem_slave_writedata -> nios2_gen2_f:jtag_debug_slave_writedata
	wire   [8:0] mm_interconnect_0_nios2_gen2_f_debug_mem_slave_address;                          // mm_interconnect_0:nios2_gen2_f_debug_mem_slave_address -> nios2_gen2_f:jtag_debug_slave_address
	wire         mm_interconnect_0_nios2_gen2_f_debug_mem_slave_write;                            // mm_interconnect_0:nios2_gen2_f_debug_mem_slave_write -> nios2_gen2_f:jtag_debug_slave_write
	wire         mm_interconnect_0_nios2_gen2_f_debug_mem_slave_read;                             // mm_interconnect_0:nios2_gen2_f_debug_mem_slave_read -> nios2_gen2_f:jtag_debug_slave_read
	wire  [31:0] mm_interconnect_0_nios2_gen2_f_debug_mem_slave_readdata;                         // nios2_gen2_f:jtag_debug_slave_readdata -> mm_interconnect_0:nios2_gen2_f_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_f_debug_mem_slave_debugaccess;                      // mm_interconnect_0:nios2_gen2_f_debug_mem_slave_debugaccess -> nios2_gen2_f:jtag_debug_slave_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_gen2_f_debug_mem_slave_byteenable;                       // mm_interconnect_0:nios2_gen2_f_debug_mem_slave_byteenable -> nios2_gen2_f:jtag_debug_slave_byteenable
	wire  [31:0] mm_interconnect_0_ipl_memory_s1_writedata;                                       // mm_interconnect_0:ipl_memory_s1_writedata -> ipl_memory:writedata
	wire  [10:0] mm_interconnect_0_ipl_memory_s1_address;                                         // mm_interconnect_0:ipl_memory_s1_address -> ipl_memory:address
	wire         mm_interconnect_0_ipl_memory_s1_chipselect;                                      // mm_interconnect_0:ipl_memory_s1_chipselect -> ipl_memory:chipselect
	wire         mm_interconnect_0_ipl_memory_s1_clken;                                           // mm_interconnect_0:ipl_memory_s1_clken -> ipl_memory:clken
	wire         mm_interconnect_0_ipl_memory_s1_write;                                           // mm_interconnect_0:ipl_memory_s1_write -> ipl_memory:write
	wire  [31:0] mm_interconnect_0_ipl_memory_s1_readdata;                                        // ipl_memory:readdata -> mm_interconnect_0:ipl_memory_s1_readdata
	wire   [3:0] mm_interconnect_0_ipl_memory_s1_byteenable;                                      // mm_interconnect_0:ipl_memory_s1_byteenable -> ipl_memory:byteenable
	wire         mm_interconnect_0_onchip_flash_0_data_waitrequest;                               // onchip_flash_0:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_0_data_waitrequest
	wire   [3:0] mm_interconnect_0_onchip_flash_0_data_burstcount;                                // mm_interconnect_0:onchip_flash_0_data_burstcount -> onchip_flash_0:avmm_data_burstcount
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_writedata;                                 // mm_interconnect_0:onchip_flash_0_data_writedata -> onchip_flash_0:avmm_data_writedata
	wire  [12:0] mm_interconnect_0_onchip_flash_0_data_address;                                   // mm_interconnect_0:onchip_flash_0_data_address -> onchip_flash_0:avmm_data_addr
	wire         mm_interconnect_0_onchip_flash_0_data_write;                                     // mm_interconnect_0:onchip_flash_0_data_write -> onchip_flash_0:avmm_data_write
	wire         mm_interconnect_0_onchip_flash_0_data_read;                                      // mm_interconnect_0:onchip_flash_0_data_read -> onchip_flash_0:avmm_data_read
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_readdata;                                  // onchip_flash_0:avmm_data_readdata -> mm_interconnect_0:onchip_flash_0_data_readdata
	wire         mm_interconnect_0_onchip_flash_0_data_readdatavalid;                             // onchip_flash_0:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_0_data_readdatavalid
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                          // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                            // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                                              // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                                           // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                                                // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                                                 // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                             // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                        // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                           // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_peripheral_bridge_s0_waitrequest;                              // peripheral_bridge:s0_waitrequest -> mm_interconnect_0:peripheral_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_0_peripheral_bridge_s0_burstcount;                               // mm_interconnect_0:peripheral_bridge_s0_burstcount -> peripheral_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_peripheral_bridge_s0_writedata;                                // mm_interconnect_0:peripheral_bridge_s0_writedata -> peripheral_bridge:s0_writedata
	wire  [15:0] mm_interconnect_0_peripheral_bridge_s0_address;                                  // mm_interconnect_0:peripheral_bridge_s0_address -> peripheral_bridge:s0_address
	wire         mm_interconnect_0_peripheral_bridge_s0_write;                                    // mm_interconnect_0:peripheral_bridge_s0_write -> peripheral_bridge:s0_write
	wire         mm_interconnect_0_peripheral_bridge_s0_read;                                     // mm_interconnect_0:peripheral_bridge_s0_read -> peripheral_bridge:s0_read
	wire  [31:0] mm_interconnect_0_peripheral_bridge_s0_readdata;                                 // peripheral_bridge:s0_readdata -> mm_interconnect_0:peripheral_bridge_s0_readdata
	wire         mm_interconnect_0_peripheral_bridge_s0_debugaccess;                              // mm_interconnect_0:peripheral_bridge_s0_debugaccess -> peripheral_bridge:s0_debugaccess
	wire         mm_interconnect_0_peripheral_bridge_s0_readdatavalid;                            // peripheral_bridge:s0_readdatavalid -> mm_interconnect_0:peripheral_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_peripheral_bridge_s0_byteenable;                               // mm_interconnect_0:peripheral_bridge_s0_byteenable -> peripheral_bridge:s0_byteenable
	wire   [0:0] peripheral_bridge_m0_burstcount;                                                 // peripheral_bridge:m0_burstcount -> mm_interconnect_1:peripheral_bridge_m0_burstcount
	wire         peripheral_bridge_m0_waitrequest;                                                // mm_interconnect_1:peripheral_bridge_m0_waitrequest -> peripheral_bridge:m0_waitrequest
	wire  [15:0] peripheral_bridge_m0_address;                                                    // peripheral_bridge:m0_address -> mm_interconnect_1:peripheral_bridge_m0_address
	wire  [31:0] peripheral_bridge_m0_writedata;                                                  // peripheral_bridge:m0_writedata -> mm_interconnect_1:peripheral_bridge_m0_writedata
	wire         peripheral_bridge_m0_write;                                                      // peripheral_bridge:m0_write -> mm_interconnect_1:peripheral_bridge_m0_write
	wire         peripheral_bridge_m0_read;                                                       // peripheral_bridge:m0_read -> mm_interconnect_1:peripheral_bridge_m0_read
	wire  [31:0] peripheral_bridge_m0_readdata;                                                   // mm_interconnect_1:peripheral_bridge_m0_readdata -> peripheral_bridge:m0_readdata
	wire         peripheral_bridge_m0_debugaccess;                                                // peripheral_bridge:m0_debugaccess -> mm_interconnect_1:peripheral_bridge_m0_debugaccess
	wire   [3:0] peripheral_bridge_m0_byteenable;                                                 // peripheral_bridge:m0_byteenable -> mm_interconnect_1:peripheral_bridge_m0_byteenable
	wire         peripheral_bridge_m0_readdatavalid;                                              // mm_interconnect_1:peripheral_bridge_m0_readdatavalid -> peripheral_bridge:m0_readdatavalid
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                                   // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                                  // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire  [15:0] mm_interconnect_1_systimer_s1_writedata;                                         // mm_interconnect_1:systimer_s1_writedata -> systimer:writedata
	wire   [2:0] mm_interconnect_1_systimer_s1_address;                                           // mm_interconnect_1:systimer_s1_address -> systimer:address
	wire         mm_interconnect_1_systimer_s1_chipselect;                                        // mm_interconnect_1:systimer_s1_chipselect -> systimer:chipselect
	wire         mm_interconnect_1_systimer_s1_write;                                             // mm_interconnect_1:systimer_s1_write -> systimer:write_n
	wire  [15:0] mm_interconnect_1_systimer_s1_readdata;                                          // systimer:readdata -> mm_interconnect_1:systimer_s1_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;                       // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;                         // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;                           // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;                        // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;                             // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;                              // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;                          // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                                              // mm_interconnect_1:led_s1_writedata -> led:writedata
	wire   [1:0] mm_interconnect_1_led_s1_address;                                                // mm_interconnect_1:led_s1_address -> led:address
	wire         mm_interconnect_1_led_s1_chipselect;                                             // mm_interconnect_1:led_s1_chipselect -> led:chipselect
	wire         mm_interconnect_1_led_s1_write;                                                  // mm_interconnect_1:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                                               // led:readdata -> mm_interconnect_1:led_s1_readdata
	wire  [31:0] mm_interconnect_1_onchip_flash_0_csr_writedata;                                  // mm_interconnect_1:onchip_flash_0_csr_writedata -> onchip_flash_0:avmm_csr_writedata
	wire   [0:0] mm_interconnect_1_onchip_flash_0_csr_address;                                    // mm_interconnect_1:onchip_flash_0_csr_address -> onchip_flash_0:avmm_csr_addr
	wire         mm_interconnect_1_onchip_flash_0_csr_write;                                      // mm_interconnect_1:onchip_flash_0_csr_write -> onchip_flash_0:avmm_csr_write
	wire         mm_interconnect_1_onchip_flash_0_csr_read;                                       // mm_interconnect_1:onchip_flash_0_csr_read -> onchip_flash_0:avmm_csr_read
	wire  [31:0] mm_interconnect_1_onchip_flash_0_csr_readdata;                                   // onchip_flash_0:avmm_csr_readdata -> mm_interconnect_1:onchip_flash_0_csr_readdata
	wire  [31:0] mm_interconnect_1_modular_adc_0_sequencer_csr_writedata;                         // mm_interconnect_1:modular_adc_0_sequencer_csr_writedata -> modular_adc_0:sequencer_csr_writedata
	wire   [0:0] mm_interconnect_1_modular_adc_0_sequencer_csr_address;                           // mm_interconnect_1:modular_adc_0_sequencer_csr_address -> modular_adc_0:sequencer_csr_address
	wire         mm_interconnect_1_modular_adc_0_sequencer_csr_write;                             // mm_interconnect_1:modular_adc_0_sequencer_csr_write -> modular_adc_0:sequencer_csr_write
	wire         mm_interconnect_1_modular_adc_0_sequencer_csr_read;                              // mm_interconnect_1:modular_adc_0_sequencer_csr_read -> modular_adc_0:sequencer_csr_read
	wire  [31:0] mm_interconnect_1_modular_adc_0_sequencer_csr_readdata;                          // modular_adc_0:sequencer_csr_readdata -> mm_interconnect_1:modular_adc_0_sequencer_csr_readdata
	wire  [31:0] mm_interconnect_1_modular_adc_0_sample_store_csr_writedata;                      // mm_interconnect_1:modular_adc_0_sample_store_csr_writedata -> modular_adc_0:sample_store_csr_writedata
	wire   [6:0] mm_interconnect_1_modular_adc_0_sample_store_csr_address;                        // mm_interconnect_1:modular_adc_0_sample_store_csr_address -> modular_adc_0:sample_store_csr_address
	wire         mm_interconnect_1_modular_adc_0_sample_store_csr_write;                          // mm_interconnect_1:modular_adc_0_sample_store_csr_write -> modular_adc_0:sample_store_csr_write
	wire         mm_interconnect_1_modular_adc_0_sample_store_csr_read;                           // mm_interconnect_1:modular_adc_0_sample_store_csr_read -> modular_adc_0:sample_store_csr_read
	wire  [31:0] mm_interconnect_1_modular_adc_0_sample_store_csr_readdata;                       // modular_adc_0:sample_store_csr_readdata -> mm_interconnect_1:modular_adc_0_sample_store_csr_readdata
	wire  [31:0] mm_interconnect_1_mmcdma_s1_writedata;                                           // mm_interconnect_1:mmcdma_s1_writedata -> mmcdma:writedata
	wire   [7:0] mm_interconnect_1_mmcdma_s1_address;                                             // mm_interconnect_1:mmcdma_s1_address -> mmcdma:address
	wire         mm_interconnect_1_mmcdma_s1_chipselect;                                          // mm_interconnect_1:mmcdma_s1_chipselect -> mmcdma:chipselect
	wire         mm_interconnect_1_mmcdma_s1_write;                                               // mm_interconnect_1:mmcdma_s1_write -> mmcdma:write
	wire         mm_interconnect_1_mmcdma_s1_read;                                                // mm_interconnect_1:mmcdma_s1_read -> mmcdma:read
	wire  [31:0] mm_interconnect_1_mmcdma_s1_readdata;                                            // mmcdma:readdata -> mm_interconnect_1:mmcdma_s1_readdata
	wire  [31:0] mm_interconnect_1_vga_s1_writedata;                                              // mm_interconnect_1:vga_s1_writedata -> vga:avs_s1_writedata
	wire   [1:0] mm_interconnect_1_vga_s1_address;                                                // mm_interconnect_1:vga_s1_address -> vga:avs_s1_address
	wire         mm_interconnect_1_vga_s1_write;                                                  // mm_interconnect_1:vga_s1_write -> vga:avs_s1_write
	wire         mm_interconnect_1_vga_s1_read;                                                   // mm_interconnect_1:vga_s1_read -> vga:avs_s1_read
	wire  [31:0] mm_interconnect_1_vga_s1_readdata;                                               // vga:avs_s1_readdata -> mm_interconnect_1:vga_s1_readdata
	wire  [31:0] nios2_gen2_f_irq_irq;                                                            // irq_mapper:sender_irq -> nios2_gen2_f:irq
	wire         irq_mapper_receiver0_irq;                                                        // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                                   // systimer:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                                        // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                               // jtag_uart:av_irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                                        // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                                               // modular_adc_0:sample_store_irq_irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver3_irq;                                                        // irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                                               // mmcdma:irq -> irq_synchronizer_003:receiver_irq
	wire         irq_mapper_receiver4_irq;                                                        // irq_synchronizer_004:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_004_receiver_irq;                                               // vga:irq_s1 -> irq_synchronizer_004:receiver_irq
	wire         rst_controller_reset_out_reset;                                                  // rst_controller:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, mm_interconnect_0:nios2_gen2_f_reset_reset_bridge_in_reset_reset, mm_interconnect_1:onchip_flash_0_nreset_reset_bridge_in_reset_reset, nios2_gen2_f:reset_n, onchip_flash_0:reset_n, rst_translator:in_reset, sdram:reset_n]
	wire         rst_controller_reset_out_reset_req;                                              // rst_controller:reset_req -> [nios2_gen2_f:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_f_debug_reset_request_reset;                                          // nios2_gen2_f:jtag_debug_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                                              // rst_controller_001:reset_out -> [ipl_memory:reset, mm_interconnect_0:ipl_memory_reset1_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                                          // rst_controller_001:reset_req -> ipl_memory:reset_req
	wire         rst_controller_002_reset_out_reset;                                              // rst_controller_002:reset_out -> [irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, jtag_uart:rst_n, led:reset_n, mm_interconnect_0:peripheral_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_1:peripheral_bridge_reset_reset_bridge_in_reset_reset, mmcdma:reset, modular_adc_0:reset_sink_reset_n, peripheral_bridge:reset, sysid:reset_n, systimer:reset_n, vga:g_reset]
	wire         rst_controller_003_reset_out_reset;                                              // rst_controller_003:reset_out -> mm_interconnect_0:vga_g_reset_reset_bridge_in_reset_reset

	testcore_nios2_gen2_f nios2_gen2_f (
		.clk                                  (clk100_clk),                                                 //                       clk.clk
		.reset_n                              (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                            (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                            (nios2_gen2_f_data_master_address),                           //               data_master.address
		.d_byteenable                         (nios2_gen2_f_data_master_byteenable),                        //                          .byteenable
		.d_read                               (nios2_gen2_f_data_master_read),                              //                          .read
		.d_readdata                           (nios2_gen2_f_data_master_readdata),                          //                          .readdata
		.d_waitrequest                        (nios2_gen2_f_data_master_waitrequest),                       //                          .waitrequest
		.d_write                              (nios2_gen2_f_data_master_write),                             //                          .write
		.d_writedata                          (nios2_gen2_f_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                      (nios2_gen2_f_data_master_readdatavalid),                     //                          .readdatavalid
		.jtag_debug_slave_debugaccess_to_roms (nios2_gen2_f_data_master_debugaccess),                       //                          .debugaccess
		.i_address                            (nios2_gen2_f_instruction_master_address),                    //        instruction_master.address
		.i_read                               (nios2_gen2_f_instruction_master_read),                       //                          .read
		.i_readdata                           (nios2_gen2_f_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                        (nios2_gen2_f_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                      (nios2_gen2_f_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                  (nios2_gen2_f_irq_irq),                                       //                       irq.irq
		.jtag_debug_resetrequest              (nios2_gen2_f_debug_reset_request_reset),                     //       debug_reset_request.reset
		.jtag_debug_slave_address             (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_address),     //           debug_mem_slave.address
		.jtag_debug_slave_byteenable          (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_byteenable),  //                          .byteenable
		.jtag_debug_slave_debugaccess         (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_debugaccess), //                          .debugaccess
		.jtag_debug_slave_read                (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_read),        //                          .read
		.jtag_debug_slave_readdata            (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_readdata),    //                          .readdata
		.jtag_debug_slave_waitrequest         (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_waitrequest), //                          .waitrequest
		.jtag_debug_slave_write               (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_write),       //                          .write
		.jtag_debug_slave_writedata           (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                      (nios2_gen2_f_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                    (nios2_gen2_f_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                         (nios2_gen2_f_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                         (nios2_gen2_f_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                         (nios2_gen2_f_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                    (nios2_gen2_f_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                     (nios2_gen2_f_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                     (nios2_gen2_f_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                 (nios2_gen2_f_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                     (nios2_gen2_f_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                     (nios2_gen2_f_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                         (nios2_gen2_f_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                    (nios2_gen2_f_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                    (nios2_gen2_f_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                     (nios2_gen2_f_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                   (nios2_gen2_f_custom_instruction_master_multi_writerc)        //                          .multi_writerc
	);

	testcore_ipl_memory ipl_memory (
		.clk        (clk100_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_ipl_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ipl_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ipl_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ipl_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ipl_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ipl_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ipl_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)      //       .reset_req
	);

	altera_onchip_flash #(
		.INIT_FILENAME               (""),
		.INIT_FILENAME_SIM           (""),
		.DEVICE_FAMILY               ("MAX 10 FPGA"),
		.PART_NAME                   ("10M08SAE144C8GES"),
		.DEVICE_ID                   ("08"),
		.SECTOR1_START_ADDR          (512),
		.SECTOR1_END_ADDR            (4607),
		.SECTOR2_START_ADDR          (4608),
		.SECTOR2_END_ADDR            (8703),
		.SECTOR3_START_ADDR          (0),
		.SECTOR3_END_ADDR            (0),
		.SECTOR4_START_ADDR          (0),
		.SECTOR4_END_ADDR            (0),
		.SECTOR5_START_ADDR          (0),
		.SECTOR5_END_ADDR            (0),
		.MIN_VALID_ADDR              (512),
		.MAX_VALID_ADDR              (8703),
		.MIN_UFM_VALID_ADDR          (512),
		.MAX_UFM_VALID_ADDR          (8703),
		.AVMM_DATA_ADDR_WIDTH        (13),
		.AVMM_DATA_BURSTCOUNT_WIDTH  (4),
		.SECTOR_READ_PROTECTION_MODE (28),
		.FLASH_SEQ_READ_DATA_COUNT   (2),
		.FLASH_ADDR_ALIGNMENT_BITS   (1),
		.FLASH_READ_CYCLE_MAX_INDEX  (3),
		.FLASH_RESET_CYCLE_MAX_INDEX (25),
		.READ_AND_WRITE_MODE         (1),
		.WRAPPING_BURST_MODE         (0),
		.IS_DUAL_BOOT                ("False")
	) onchip_flash_0 (
		.clock                   (clk100_clk),                                          //    clk.clk
		.reset_n                 (~rst_controller_reset_out_reset),                     // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_onchip_flash_0_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_onchip_flash_0_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_0_onchip_flash_0_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_0_onchip_flash_0_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_0_onchip_flash_0_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_onchip_flash_0_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_onchip_flash_0_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_onchip_flash_0_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_1_onchip_flash_0_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_1_onchip_flash_0_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_1_onchip_flash_0_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_1_onchip_flash_0_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_1_onchip_flash_0_csr_readdata)        //       .readdata
	);

	testcore_sysid sysid (
		.clock    (clk40_clk),                                      //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	testcore_systimer systimer (
		.clk        (clk40_clk),                                //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.address    (mm_interconnect_1_systimer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_systimer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_systimer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_systimer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_systimer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)             //   irq.irq
	);

	testcore_jtag_uart jtag_uart (
		.clk            (clk40_clk),                                                 //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_001_receiver_irq)                          //               irq.irq
	);

	testcore_led led (
		.clk        (clk40_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (16),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) peripheral_bridge (
		.clk              (clk40_clk),                                            //   clk.clk
		.reset            (rst_controller_002_reset_out_reset),                   // reset.reset
		.s0_waitrequest   (mm_interconnect_0_peripheral_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_peripheral_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_peripheral_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_peripheral_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_peripheral_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_peripheral_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_peripheral_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_peripheral_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_peripheral_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_peripheral_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (peripheral_bridge_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (peripheral_bridge_m0_readdata),                        //      .readdata
		.m0_readdatavalid (peripheral_bridge_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (peripheral_bridge_m0_burstcount),                      //      .burstcount
		.m0_writedata     (peripheral_bridge_m0_writedata),                       //      .writedata
		.m0_address       (peripheral_bridge_m0_address),                         //      .address
		.m0_write         (peripheral_bridge_m0_write),                           //      .write
		.m0_read          (peripheral_bridge_m0_read),                            //      .read
		.m0_byteenable    (peripheral_bridge_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (peripheral_bridge_m0_debugaccess)                      //      .debugaccess
	);

	testcore_sdram sdram (
		.clk            (clk100_clk),                               //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdr_addr),                                 //  wire.export
		.zs_ba          (sdr_ba),                                   //      .export
		.zs_cas_n       (sdr_cas_n),                                //      .export
		.zs_cke         (sdr_cke),                                  //      .export
		.zs_cs_n        (sdr_cs_n),                                 //      .export
		.zs_dq          (sdr_dq),                                   //      .export
		.zs_dqm         (sdr_dqm),                                  //      .export
		.zs_ras_n       (sdr_ras_n),                                //      .export
		.zs_we_n        (sdr_we_n)                                  //      .export
	);

	testcore_modular_adc_0 modular_adc_0 (
		.clock_clk                  (clk40_clk),                                                  //            clock.clk
		.reset_sink_reset_n         (~rst_controller_002_reset_out_reset),                        //       reset_sink.reset_n
		.adc_pll_clock_clk          (clk40_clk),                                                  //    adc_pll_clock.clk
		.adc_pll_locked_export      (adc_pll_locked_export),                                      //   adc_pll_locked.export
		.sequencer_csr_address      (mm_interconnect_1_modular_adc_0_sequencer_csr_address),      //    sequencer_csr.address
		.sequencer_csr_read         (mm_interconnect_1_modular_adc_0_sequencer_csr_read),         //                 .read
		.sequencer_csr_write        (mm_interconnect_1_modular_adc_0_sequencer_csr_write),        //                 .write
		.sequencer_csr_writedata    (mm_interconnect_1_modular_adc_0_sequencer_csr_writedata),    //                 .writedata
		.sequencer_csr_readdata     (mm_interconnect_1_modular_adc_0_sequencer_csr_readdata),     //                 .readdata
		.sample_store_csr_address   (mm_interconnect_1_modular_adc_0_sample_store_csr_address),   // sample_store_csr.address
		.sample_store_csr_read      (mm_interconnect_1_modular_adc_0_sample_store_csr_read),      //                 .read
		.sample_store_csr_write     (mm_interconnect_1_modular_adc_0_sample_store_csr_write),     //                 .write
		.sample_store_csr_writedata (mm_interconnect_1_modular_adc_0_sample_store_csr_writedata), //                 .writedata
		.sample_store_csr_readdata  (mm_interconnect_1_modular_adc_0_sample_store_csr_readdata),  //                 .readdata
		.sample_store_irq_irq       (irq_synchronizer_002_receiver_irq)                           // sample_store_irq.irq
	);

	pixelsimd pixelsimd (
		.dataa  (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave_0.dataa
		.datab  (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //                                .datab
		.result (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_result), //                                .result
		.clk    (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //                                .clk
		.clk_en (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //                                .clk_en
		.reset  (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //                                .reset
		.start  (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_start),  //                                .start
		.done   (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_done),   //                                .done
		.n      (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_n)       //                                .n
	);

	avalonif_mmcdma #(
		.SYSTEMCLOCKINFO (40000000)
	) mmcdma (
		.clk        (clk40_clk),                              //       clock_reset.clk
		.reset      (rst_controller_002_reset_out_reset),     // clock_reset_reset.reset
		.chipselect (mm_interconnect_1_mmcdma_s1_chipselect), //                s1.chipselect
		.address    (mm_interconnect_1_mmcdma_s1_address),    //                  .address
		.read       (mm_interconnect_1_mmcdma_s1_read),       //                  .read
		.readdata   (mm_interconnect_1_mmcdma_s1_readdata),   //                  .readdata
		.write      (mm_interconnect_1_mmcdma_s1_write),      //                  .write
		.writedata  (mm_interconnect_1_mmcdma_s1_writedata),  //                  .writedata
		.MMC_nCS    (mmc_nCS),                                //       conduit_end.export
		.MMC_SCK    (mmc_SCK),                                //                  .export
		.MMC_SDO    (mmc_SDO),                                //                  .export
		.MMC_SDI    (mmc_SDI),                                //                  .export
		.MMC_CD     (mmc_CD),                                 //                  .export
		.MMC_WP     (mmc_WP),                                 //                  .export
		.irq        (irq_synchronizer_003_receiver_irq)       //  interrupt_sender.irq
	);

	vga_component #(
		.LINEOFFSETBYTES (2048),
		.H_TOTAL         (794),
		.H_SYNC          (96),
		.H_BACKP         (48),
		.H_ACTIVE        (640),
		.V_TOTAL         (525),
		.V_SYNC          (2),
		.V_BACKP         (33),
		.V_ACTIVE        (480)
	) vga (
		.video_clk            (vga_clk),                            //     ext.export
		.video_rout           (vga_rout),                           //        .export
		.video_gout           (vga_gout),                           //        .export
		.video_bout           (vga_bout),                           //        .export
		.video_hsync_n        (vga_hsync_n),                        //        .export
		.video_vsync_n        (vga_vsync_n),                        //        .export
		.video_enable         (vga_enable),                         //        .export
		.avm_m1_address       (vga_m1_address),                     //      m1.address
		.avm_m1_waitrequest   (vga_m1_waitrequest),                 //        .waitrequest
		.avm_m1_burstcount    (vga_m1_burstcount),                  //        .burstcount
		.avm_m1_read          (vga_m1_read),                        //        .read
		.avm_m1_readdata      (vga_m1_readdata),                    //        .readdata
		.avm_m1_readdatavalid (vga_m1_readdatavalid),               //        .readdatavalid
		.avs_s1_address       (mm_interconnect_1_vga_s1_address),   //      s1.address
		.avs_s1_read          (mm_interconnect_1_vga_s1_read),      //        .read
		.avs_s1_readdata      (mm_interconnect_1_vga_s1_readdata),  //        .readdata
		.avs_s1_write         (mm_interconnect_1_vga_s1_write),     //        .write
		.avs_s1_writedata     (mm_interconnect_1_vga_s1_writedata), //        .writedata
		.irq_s1               (irq_synchronizer_004_receiver_irq),  //     irq.irq
		.s1_clk               (clk40_clk),                          //   s_clk.clk
		.m1_clk               (clk100_clk),                         //   m_clk.clk
		.g_reset              (rst_controller_002_reset_out_reset)  // g_reset.reset
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_gen2_f_custom_instruction_master_translator (
		.ci_slave_result           (),                                                                            //        ci_slave.result
		.ci_slave_multi_clk        (nios2_gen2_f_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_gen2_f_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_gen2_f_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_gen2_f_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_gen2_f_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_gen2_f_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios2_gen2_f_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios2_gen2_f_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios2_gen2_f_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios2_gen2_f_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios2_gen2_f_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios2_gen2_f_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios2_gen2_f_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios2_gen2_f_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios2_gen2_f_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios2_gen2_f_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_result     (),                                                                            //  comb_ci_master.result
		.multi_ci_master_clk       (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_dataa            (32'b00000000000000000000000000000000),                                        //     (terminated)
		.ci_slave_datab            (32'b00000000000000000000000000000000),                                        //     (terminated)
		.ci_slave_n                (8'b00000000),                                                                 //     (terminated)
		.ci_slave_readra           (1'b0),                                                                        //     (terminated)
		.ci_slave_readrb           (1'b0),                                                                        //     (terminated)
		.ci_slave_writerc          (1'b0),                                                                        //     (terminated)
		.ci_slave_a                (5'b00000),                                                                    //     (terminated)
		.ci_slave_b                (5'b00000),                                                                    //     (terminated)
		.ci_slave_c                (5'b00000),                                                                    //     (terminated)
		.ci_slave_ipending         (32'b00000000000000000000000000000000),                                        //     (terminated)
		.ci_slave_estatus          (1'b0),                                                                        //     (terminated)
		.comb_ci_master_dataa      (),                                                                            //     (terminated)
		.comb_ci_master_datab      (),                                                                            //     (terminated)
		.comb_ci_master_n          (),                                                                            //     (terminated)
		.comb_ci_master_readra     (),                                                                            //     (terminated)
		.comb_ci_master_readrb     (),                                                                            //     (terminated)
		.comb_ci_master_writerc    (),                                                                            //     (terminated)
		.comb_ci_master_a          (),                                                                            //     (terminated)
		.comb_ci_master_b          (),                                                                            //     (terminated)
		.comb_ci_master_c          (),                                                                            //     (terminated)
		.comb_ci_master_ipending   (),                                                                            //     (terminated)
		.comb_ci_master_estatus    ()                                                                             //     (terminated)
	);

	testcore_nios2_gen2_f_custom_instruction_master_multi_xconnect nios2_gen2_f_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                            //           .ipending
		.ci_slave_estatus     (),                                                                            //           .estatus
		.ci_slave_clk         (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_gen2_f_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_gen2_f_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios2_gen2_f_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_n),      //          .n
		.ci_master_clk       (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios2_gen2_f_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_readra    (),                                                                                // (terminated)
		.ci_master_readrb    (),                                                                                // (terminated)
		.ci_master_writerc   (),                                                                                // (terminated)
		.ci_master_a         (),                                                                                // (terminated)
		.ci_master_b         (),                                                                                // (terminated)
		.ci_master_c         (),                                                                                // (terminated)
		.ci_master_ipending  (),                                                                                // (terminated)
		.ci_master_estatus   (),                                                                                // (terminated)
		.ci_master_reset_req ()                                                                                 // (terminated)
	);

	testcore_mm_interconnect_0 mm_interconnect_0 (
		.clk_core_clk_clk                                    (clk100_clk),                                                 //                                  clk_core_clk.clk
		.clk_peri_clk_clk                                    (clk40_clk),                                                  //                                  clk_peri_clk.clk
		.ipl_memory_reset1_reset_bridge_in_reset_reset       (rst_controller_001_reset_out_reset),                         //       ipl_memory_reset1_reset_bridge_in_reset.reset
		.nios2_gen2_f_reset_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                             //      nios2_gen2_f_reset_reset_bridge_in_reset.reset
		.peripheral_bridge_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                         // peripheral_bridge_reset_reset_bridge_in_reset.reset
		.vga_g_reset_reset_bridge_in_reset_reset             (rst_controller_003_reset_out_reset),                         //             vga_g_reset_reset_bridge_in_reset.reset
		.nios2_gen2_f_data_master_address                    (nios2_gen2_f_data_master_address),                           //                      nios2_gen2_f_data_master.address
		.nios2_gen2_f_data_master_waitrequest                (nios2_gen2_f_data_master_waitrequest),                       //                                              .waitrequest
		.nios2_gen2_f_data_master_byteenable                 (nios2_gen2_f_data_master_byteenable),                        //                                              .byteenable
		.nios2_gen2_f_data_master_read                       (nios2_gen2_f_data_master_read),                              //                                              .read
		.nios2_gen2_f_data_master_readdata                   (nios2_gen2_f_data_master_readdata),                          //                                              .readdata
		.nios2_gen2_f_data_master_readdatavalid              (nios2_gen2_f_data_master_readdatavalid),                     //                                              .readdatavalid
		.nios2_gen2_f_data_master_write                      (nios2_gen2_f_data_master_write),                             //                                              .write
		.nios2_gen2_f_data_master_writedata                  (nios2_gen2_f_data_master_writedata),                         //                                              .writedata
		.nios2_gen2_f_data_master_debugaccess                (nios2_gen2_f_data_master_debugaccess),                       //                                              .debugaccess
		.nios2_gen2_f_instruction_master_address             (nios2_gen2_f_instruction_master_address),                    //               nios2_gen2_f_instruction_master.address
		.nios2_gen2_f_instruction_master_waitrequest         (nios2_gen2_f_instruction_master_waitrequest),                //                                              .waitrequest
		.nios2_gen2_f_instruction_master_read                (nios2_gen2_f_instruction_master_read),                       //                                              .read
		.nios2_gen2_f_instruction_master_readdata            (nios2_gen2_f_instruction_master_readdata),                   //                                              .readdata
		.nios2_gen2_f_instruction_master_readdatavalid       (nios2_gen2_f_instruction_master_readdatavalid),              //                                              .readdatavalid
		.vga_m1_address                                      (vga_m1_address),                                             //                                        vga_m1.address
		.vga_m1_waitrequest                                  (vga_m1_waitrequest),                                         //                                              .waitrequest
		.vga_m1_burstcount                                   (vga_m1_burstcount),                                          //                                              .burstcount
		.vga_m1_read                                         (vga_m1_read),                                                //                                              .read
		.vga_m1_readdata                                     (vga_m1_readdata),                                            //                                              .readdata
		.vga_m1_readdatavalid                                (vga_m1_readdatavalid),                                       //                                              .readdatavalid
		.ipl_memory_s1_address                               (mm_interconnect_0_ipl_memory_s1_address),                    //                                 ipl_memory_s1.address
		.ipl_memory_s1_write                                 (mm_interconnect_0_ipl_memory_s1_write),                      //                                              .write
		.ipl_memory_s1_readdata                              (mm_interconnect_0_ipl_memory_s1_readdata),                   //                                              .readdata
		.ipl_memory_s1_writedata                             (mm_interconnect_0_ipl_memory_s1_writedata),                  //                                              .writedata
		.ipl_memory_s1_byteenable                            (mm_interconnect_0_ipl_memory_s1_byteenable),                 //                                              .byteenable
		.ipl_memory_s1_chipselect                            (mm_interconnect_0_ipl_memory_s1_chipselect),                 //                                              .chipselect
		.ipl_memory_s1_clken                                 (mm_interconnect_0_ipl_memory_s1_clken),                      //                                              .clken
		.nios2_gen2_f_debug_mem_slave_address                (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_address),     //                  nios2_gen2_f_debug_mem_slave.address
		.nios2_gen2_f_debug_mem_slave_write                  (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_write),       //                                              .write
		.nios2_gen2_f_debug_mem_slave_read                   (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_read),        //                                              .read
		.nios2_gen2_f_debug_mem_slave_readdata               (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_readdata),    //                                              .readdata
		.nios2_gen2_f_debug_mem_slave_writedata              (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_writedata),   //                                              .writedata
		.nios2_gen2_f_debug_mem_slave_byteenable             (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_byteenable),  //                                              .byteenable
		.nios2_gen2_f_debug_mem_slave_waitrequest            (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_waitrequest), //                                              .waitrequest
		.nios2_gen2_f_debug_mem_slave_debugaccess            (mm_interconnect_0_nios2_gen2_f_debug_mem_slave_debugaccess), //                                              .debugaccess
		.onchip_flash_0_data_address                         (mm_interconnect_0_onchip_flash_0_data_address),              //                           onchip_flash_0_data.address
		.onchip_flash_0_data_write                           (mm_interconnect_0_onchip_flash_0_data_write),                //                                              .write
		.onchip_flash_0_data_read                            (mm_interconnect_0_onchip_flash_0_data_read),                 //                                              .read
		.onchip_flash_0_data_readdata                        (mm_interconnect_0_onchip_flash_0_data_readdata),             //                                              .readdata
		.onchip_flash_0_data_writedata                       (mm_interconnect_0_onchip_flash_0_data_writedata),            //                                              .writedata
		.onchip_flash_0_data_burstcount                      (mm_interconnect_0_onchip_flash_0_data_burstcount),           //                                              .burstcount
		.onchip_flash_0_data_readdatavalid                   (mm_interconnect_0_onchip_flash_0_data_readdatavalid),        //                                              .readdatavalid
		.onchip_flash_0_data_waitrequest                     (mm_interconnect_0_onchip_flash_0_data_waitrequest),          //                                              .waitrequest
		.peripheral_bridge_s0_address                        (mm_interconnect_0_peripheral_bridge_s0_address),             //                          peripheral_bridge_s0.address
		.peripheral_bridge_s0_write                          (mm_interconnect_0_peripheral_bridge_s0_write),               //                                              .write
		.peripheral_bridge_s0_read                           (mm_interconnect_0_peripheral_bridge_s0_read),                //                                              .read
		.peripheral_bridge_s0_readdata                       (mm_interconnect_0_peripheral_bridge_s0_readdata),            //                                              .readdata
		.peripheral_bridge_s0_writedata                      (mm_interconnect_0_peripheral_bridge_s0_writedata),           //                                              .writedata
		.peripheral_bridge_s0_burstcount                     (mm_interconnect_0_peripheral_bridge_s0_burstcount),          //                                              .burstcount
		.peripheral_bridge_s0_byteenable                     (mm_interconnect_0_peripheral_bridge_s0_byteenable),          //                                              .byteenable
		.peripheral_bridge_s0_readdatavalid                  (mm_interconnect_0_peripheral_bridge_s0_readdatavalid),       //                                              .readdatavalid
		.peripheral_bridge_s0_waitrequest                    (mm_interconnect_0_peripheral_bridge_s0_waitrequest),         //                                              .waitrequest
		.peripheral_bridge_s0_debugaccess                    (mm_interconnect_0_peripheral_bridge_s0_debugaccess),         //                                              .debugaccess
		.sdram_s1_address                                    (mm_interconnect_0_sdram_s1_address),                         //                                      sdram_s1.address
		.sdram_s1_write                                      (mm_interconnect_0_sdram_s1_write),                           //                                              .write
		.sdram_s1_read                                       (mm_interconnect_0_sdram_s1_read),                            //                                              .read
		.sdram_s1_readdata                                   (mm_interconnect_0_sdram_s1_readdata),                        //                                              .readdata
		.sdram_s1_writedata                                  (mm_interconnect_0_sdram_s1_writedata),                       //                                              .writedata
		.sdram_s1_byteenable                                 (mm_interconnect_0_sdram_s1_byteenable),                      //                                              .byteenable
		.sdram_s1_readdatavalid                              (mm_interconnect_0_sdram_s1_readdatavalid),                   //                                              .readdatavalid
		.sdram_s1_waitrequest                                (mm_interconnect_0_sdram_s1_waitrequest),                     //                                              .waitrequest
		.sdram_s1_chipselect                                 (mm_interconnect_0_sdram_s1_chipselect)                       //                                              .chipselect
	);

	testcore_mm_interconnect_1 mm_interconnect_1 (
		.clk_core_clk_clk                                    (clk100_clk),                                                 //                                  clk_core_clk.clk
		.clk_peri_clk_clk                                    (clk40_clk),                                                  //                                  clk_peri_clk.clk
		.onchip_flash_0_nreset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                             //   onchip_flash_0_nreset_reset_bridge_in_reset.reset
		.peripheral_bridge_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                         // peripheral_bridge_reset_reset_bridge_in_reset.reset
		.peripheral_bridge_m0_address                        (peripheral_bridge_m0_address),                               //                          peripheral_bridge_m0.address
		.peripheral_bridge_m0_waitrequest                    (peripheral_bridge_m0_waitrequest),                           //                                              .waitrequest
		.peripheral_bridge_m0_burstcount                     (peripheral_bridge_m0_burstcount),                            //                                              .burstcount
		.peripheral_bridge_m0_byteenable                     (peripheral_bridge_m0_byteenable),                            //                                              .byteenable
		.peripheral_bridge_m0_read                           (peripheral_bridge_m0_read),                                  //                                              .read
		.peripheral_bridge_m0_readdata                       (peripheral_bridge_m0_readdata),                              //                                              .readdata
		.peripheral_bridge_m0_readdatavalid                  (peripheral_bridge_m0_readdatavalid),                         //                                              .readdatavalid
		.peripheral_bridge_m0_write                          (peripheral_bridge_m0_write),                                 //                                              .write
		.peripheral_bridge_m0_writedata                      (peripheral_bridge_m0_writedata),                             //                                              .writedata
		.peripheral_bridge_m0_debugaccess                    (peripheral_bridge_m0_debugaccess),                           //                                              .debugaccess
		.jtag_uart_avalon_jtag_slave_address                 (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),      //                   jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),        //                                              .write
		.jtag_uart_avalon_jtag_slave_read                    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),         //                                              .read
		.jtag_uart_avalon_jtag_slave_readdata                (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),     //                                              .readdata
		.jtag_uart_avalon_jtag_slave_writedata               (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),    //                                              .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest             (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest),  //                                              .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect              (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),   //                                              .chipselect
		.led_s1_address                                      (mm_interconnect_1_led_s1_address),                           //                                        led_s1.address
		.led_s1_write                                        (mm_interconnect_1_led_s1_write),                             //                                              .write
		.led_s1_readdata                                     (mm_interconnect_1_led_s1_readdata),                          //                                              .readdata
		.led_s1_writedata                                    (mm_interconnect_1_led_s1_writedata),                         //                                              .writedata
		.led_s1_chipselect                                   (mm_interconnect_1_led_s1_chipselect),                        //                                              .chipselect
		.mmcdma_s1_address                                   (mm_interconnect_1_mmcdma_s1_address),                        //                                     mmcdma_s1.address
		.mmcdma_s1_write                                     (mm_interconnect_1_mmcdma_s1_write),                          //                                              .write
		.mmcdma_s1_read                                      (mm_interconnect_1_mmcdma_s1_read),                           //                                              .read
		.mmcdma_s1_readdata                                  (mm_interconnect_1_mmcdma_s1_readdata),                       //                                              .readdata
		.mmcdma_s1_writedata                                 (mm_interconnect_1_mmcdma_s1_writedata),                      //                                              .writedata
		.mmcdma_s1_chipselect                                (mm_interconnect_1_mmcdma_s1_chipselect),                     //                                              .chipselect
		.modular_adc_0_sample_store_csr_address              (mm_interconnect_1_modular_adc_0_sample_store_csr_address),   //                modular_adc_0_sample_store_csr.address
		.modular_adc_0_sample_store_csr_write                (mm_interconnect_1_modular_adc_0_sample_store_csr_write),     //                                              .write
		.modular_adc_0_sample_store_csr_read                 (mm_interconnect_1_modular_adc_0_sample_store_csr_read),      //                                              .read
		.modular_adc_0_sample_store_csr_readdata             (mm_interconnect_1_modular_adc_0_sample_store_csr_readdata),  //                                              .readdata
		.modular_adc_0_sample_store_csr_writedata            (mm_interconnect_1_modular_adc_0_sample_store_csr_writedata), //                                              .writedata
		.modular_adc_0_sequencer_csr_address                 (mm_interconnect_1_modular_adc_0_sequencer_csr_address),      //                   modular_adc_0_sequencer_csr.address
		.modular_adc_0_sequencer_csr_write                   (mm_interconnect_1_modular_adc_0_sequencer_csr_write),        //                                              .write
		.modular_adc_0_sequencer_csr_read                    (mm_interconnect_1_modular_adc_0_sequencer_csr_read),         //                                              .read
		.modular_adc_0_sequencer_csr_readdata                (mm_interconnect_1_modular_adc_0_sequencer_csr_readdata),     //                                              .readdata
		.modular_adc_0_sequencer_csr_writedata               (mm_interconnect_1_modular_adc_0_sequencer_csr_writedata),    //                                              .writedata
		.onchip_flash_0_csr_address                          (mm_interconnect_1_onchip_flash_0_csr_address),               //                            onchip_flash_0_csr.address
		.onchip_flash_0_csr_write                            (mm_interconnect_1_onchip_flash_0_csr_write),                 //                                              .write
		.onchip_flash_0_csr_read                             (mm_interconnect_1_onchip_flash_0_csr_read),                  //                                              .read
		.onchip_flash_0_csr_readdata                         (mm_interconnect_1_onchip_flash_0_csr_readdata),              //                                              .readdata
		.onchip_flash_0_csr_writedata                        (mm_interconnect_1_onchip_flash_0_csr_writedata),             //                                              .writedata
		.sysid_control_slave_address                         (mm_interconnect_1_sysid_control_slave_address),              //                           sysid_control_slave.address
		.sysid_control_slave_readdata                        (mm_interconnect_1_sysid_control_slave_readdata),             //                                              .readdata
		.systimer_s1_address                                 (mm_interconnect_1_systimer_s1_address),                      //                                   systimer_s1.address
		.systimer_s1_write                                   (mm_interconnect_1_systimer_s1_write),                        //                                              .write
		.systimer_s1_readdata                                (mm_interconnect_1_systimer_s1_readdata),                     //                                              .readdata
		.systimer_s1_writedata                               (mm_interconnect_1_systimer_s1_writedata),                    //                                              .writedata
		.systimer_s1_chipselect                              (mm_interconnect_1_systimer_s1_chipselect),                   //                                              .chipselect
		.vga_s1_address                                      (mm_interconnect_1_vga_s1_address),                           //                                        vga_s1.address
		.vga_s1_write                                        (mm_interconnect_1_vga_s1_write),                             //                                              .write
		.vga_s1_read                                         (mm_interconnect_1_vga_s1_read),                              //                                              .read
		.vga_s1_readdata                                     (mm_interconnect_1_vga_s1_readdata),                          //                                              .readdata
		.vga_s1_writedata                                    (mm_interconnect_1_vga_s1_writedata)                          //                                              .writedata
	);

	testcore_irq_mapper irq_mapper (
		.clk           (clk100_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (nios2_gen2_f_irq_irq)            //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk40_clk),                          //       receiver_clk.clk
		.sender_clk     (clk100_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk40_clk),                          //       receiver_clk.clk
		.sender_clk     (clk100_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk40_clk),                          //       receiver_clk.clk
		.sender_clk     (clk100_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk40_clk),                          //       receiver_clk.clk
		.sender_clk     (clk100_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (clk40_clk),                          //       receiver_clk.clk
		.sender_clk     (clk100_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_f_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk100_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk100_clk),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk40_clk),                          //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk100_clk),                         //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
