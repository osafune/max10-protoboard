// testcore.v

// Generated using ACDS version 14.0 209 at 2014.11.14.01:06:16

`timescale 1 ps / 1 ps
module testcore (
		input  wire        clk100_clk,            //         clk100.clk
		input  wire        reset_reset_n,         //          reset.reset_n
		output wire        led_export,            //            led.export
		inout  wire [27:0] gpio_export,           //           gpio.export
		input  wire        clk40_clk,             //          clk40.clk
		output wire [12:0] sdr_addr,              //            sdr.addr
		output wire [1:0]  sdr_ba,                //               .ba
		output wire        sdr_cas_n,             //               .cas_n
		output wire        sdr_cke,               //               .cke
		output wire        sdr_cs_n,              //               .cs_n
		inout  wire [15:0] sdr_dq,                //               .dq
		output wire [1:0]  sdr_dqm,               //               .dqm
		output wire        sdr_ras_n,             //               .ras_n
		output wire        sdr_we_n,              //               .we_n
		input  wire        adc_pll_locked_export  // adc_pll_locked.export
	);

	wire         nios2_gen2_0_instruction_master_waitrequest;                // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [27:0] nios2_gen2_0_instruction_master_address;                    // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                       // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_readdatavalid;              // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         nios2_gen2_0_data_master_waitrequest;                       // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire  [31:0] nios2_gen2_0_data_master_writedata;                         // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [28:0] nios2_gen2_0_data_master_address;                           // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire         nios2_gen2_0_data_master_write;                             // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire         nios2_gen2_0_data_master_read;                              // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire  [31:0] nios2_gen2_0_data_master_readdata;                          // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_debugaccess;                       // nios2_gen2_0:jtag_debug_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire         nios2_gen2_0_data_master_readdatavalid;                     // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                        // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest; // nios2_gen2_0:jtag_debug_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:jtag_debug_slave_writedata
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:jtag_debug_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:jtag_debug_slave_write
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:jtag_debug_slave_read
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;    // nios2_gen2_0:jtag_debug_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:jtag_debug_slave_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:jtag_debug_slave_byteenable
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;            // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire  [11:0] mm_interconnect_0_onchip_memory2_0_s1_address;              // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;           // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;             // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;           // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_flash_0_data_waitrequest;          // onchip_flash_0:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_0_data_waitrequest
	wire   [3:0] mm_interconnect_0_onchip_flash_0_data_burstcount;           // mm_interconnect_0:onchip_flash_0_data_burstcount -> onchip_flash_0:avmm_data_burstcount
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_writedata;            // mm_interconnect_0:onchip_flash_0_data_writedata -> onchip_flash_0:avmm_data_writedata
	wire  [12:0] mm_interconnect_0_onchip_flash_0_data_address;              // mm_interconnect_0:onchip_flash_0_data_address -> onchip_flash_0:avmm_data_addr
	wire         mm_interconnect_0_onchip_flash_0_data_write;                // mm_interconnect_0:onchip_flash_0_data_write -> onchip_flash_0:avmm_data_write
	wire         mm_interconnect_0_onchip_flash_0_data_read;                 // mm_interconnect_0:onchip_flash_0_data_read -> onchip_flash_0:avmm_data_read
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_readdata;             // onchip_flash_0:avmm_data_readdata -> mm_interconnect_0:onchip_flash_0_data_readdata
	wire         mm_interconnect_0_onchip_flash_0_data_readdatavalid;        // onchip_flash_0:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_0_data_readdatavalid
	wire         mm_interconnect_0_sdram_s1_waitrequest;                     // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                       // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                         // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                      // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                           // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                            // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                        // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                   // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                      // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_peripheral_bridge_s0_waitrequest;         // peripheral_bridge:s0_waitrequest -> mm_interconnect_0:peripheral_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_0_peripheral_bridge_s0_burstcount;          // mm_interconnect_0:peripheral_bridge_s0_burstcount -> peripheral_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_peripheral_bridge_s0_writedata;           // mm_interconnect_0:peripheral_bridge_s0_writedata -> peripheral_bridge:s0_writedata
	wire  [15:0] mm_interconnect_0_peripheral_bridge_s0_address;             // mm_interconnect_0:peripheral_bridge_s0_address -> peripheral_bridge:s0_address
	wire         mm_interconnect_0_peripheral_bridge_s0_write;               // mm_interconnect_0:peripheral_bridge_s0_write -> peripheral_bridge:s0_write
	wire         mm_interconnect_0_peripheral_bridge_s0_read;                // mm_interconnect_0:peripheral_bridge_s0_read -> peripheral_bridge:s0_read
	wire  [31:0] mm_interconnect_0_peripheral_bridge_s0_readdata;            // peripheral_bridge:s0_readdata -> mm_interconnect_0:peripheral_bridge_s0_readdata
	wire         mm_interconnect_0_peripheral_bridge_s0_debugaccess;         // mm_interconnect_0:peripheral_bridge_s0_debugaccess -> peripheral_bridge:s0_debugaccess
	wire         mm_interconnect_0_peripheral_bridge_s0_readdatavalid;       // peripheral_bridge:s0_readdatavalid -> mm_interconnect_0:peripheral_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_peripheral_bridge_s0_byteenable;          // mm_interconnect_0:peripheral_bridge_s0_byteenable -> peripheral_bridge:s0_byteenable
	wire   [0:0] peripheral_bridge_m0_burstcount;                            // peripheral_bridge:m0_burstcount -> mm_interconnect_1:peripheral_bridge_m0_burstcount
	wire         peripheral_bridge_m0_waitrequest;                           // mm_interconnect_1:peripheral_bridge_m0_waitrequest -> peripheral_bridge:m0_waitrequest
	wire  [15:0] peripheral_bridge_m0_address;                               // peripheral_bridge:m0_address -> mm_interconnect_1:peripheral_bridge_m0_address
	wire  [31:0] peripheral_bridge_m0_writedata;                             // peripheral_bridge:m0_writedata -> mm_interconnect_1:peripheral_bridge_m0_writedata
	wire         peripheral_bridge_m0_write;                                 // peripheral_bridge:m0_write -> mm_interconnect_1:peripheral_bridge_m0_write
	wire         peripheral_bridge_m0_read;                                  // peripheral_bridge:m0_read -> mm_interconnect_1:peripheral_bridge_m0_read
	wire  [31:0] peripheral_bridge_m0_readdata;                              // mm_interconnect_1:peripheral_bridge_m0_readdata -> peripheral_bridge:m0_readdata
	wire         peripheral_bridge_m0_debugaccess;                           // peripheral_bridge:m0_debugaccess -> mm_interconnect_1:peripheral_bridge_m0_debugaccess
	wire   [3:0] peripheral_bridge_m0_byteenable;                            // peripheral_bridge:m0_byteenable -> mm_interconnect_1:peripheral_bridge_m0_byteenable
	wire         peripheral_bridge_m0_readdatavalid;                         // mm_interconnect_1:peripheral_bridge_m0_readdatavalid -> peripheral_bridge:m0_readdatavalid
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;              // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;             // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire  [15:0] mm_interconnect_1_systimer_s1_writedata;                    // mm_interconnect_1:systimer_s1_writedata -> systimer:writedata
	wire   [2:0] mm_interconnect_1_systimer_s1_address;                      // mm_interconnect_1:systimer_s1_address -> systimer:address
	wire         mm_interconnect_1_systimer_s1_chipselect;                   // mm_interconnect_1:systimer_s1_chipselect -> systimer:chipselect
	wire         mm_interconnect_1_systimer_s1_write;                        // mm_interconnect_1:systimer_s1_write -> systimer:write_n
	wire  [15:0] mm_interconnect_1_systimer_s1_readdata;                     // systimer:readdata -> mm_interconnect_1:systimer_s1_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;  // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;    // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;      // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;   // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;        // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;         // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;     // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                         // mm_interconnect_1:led_s1_writedata -> led:writedata
	wire   [1:0] mm_interconnect_1_led_s1_address;                           // mm_interconnect_1:led_s1_address -> led:address
	wire         mm_interconnect_1_led_s1_chipselect;                        // mm_interconnect_1:led_s1_chipselect -> led:chipselect
	wire         mm_interconnect_1_led_s1_write;                             // mm_interconnect_1:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                          // led:readdata -> mm_interconnect_1:led_s1_readdata
	wire  [31:0] mm_interconnect_1_gpio_s1_writedata;                        // mm_interconnect_1:gpio_s1_writedata -> gpio:writedata
	wire   [1:0] mm_interconnect_1_gpio_s1_address;                          // mm_interconnect_1:gpio_s1_address -> gpio:address
	wire         mm_interconnect_1_gpio_s1_chipselect;                       // mm_interconnect_1:gpio_s1_chipselect -> gpio:chipselect
	wire         mm_interconnect_1_gpio_s1_write;                            // mm_interconnect_1:gpio_s1_write -> gpio:write_n
	wire  [31:0] mm_interconnect_1_gpio_s1_readdata;                         // gpio:readdata -> mm_interconnect_1:gpio_s1_readdata
	wire  [31:0] mm_interconnect_1_onchip_flash_0_csr_writedata;             // mm_interconnect_1:onchip_flash_0_csr_writedata -> onchip_flash_0:avmm_csr_writedata
	wire   [0:0] mm_interconnect_1_onchip_flash_0_csr_address;               // mm_interconnect_1:onchip_flash_0_csr_address -> onchip_flash_0:avmm_csr_addr
	wire         mm_interconnect_1_onchip_flash_0_csr_write;                 // mm_interconnect_1:onchip_flash_0_csr_write -> onchip_flash_0:avmm_csr_write
	wire         mm_interconnect_1_onchip_flash_0_csr_read;                  // mm_interconnect_1:onchip_flash_0_csr_read -> onchip_flash_0:avmm_csr_read
	wire  [31:0] mm_interconnect_1_onchip_flash_0_csr_readdata;              // onchip_flash_0:avmm_csr_readdata -> mm_interconnect_1:onchip_flash_0_csr_readdata
	wire  [31:0] mm_interconnect_1_modular_adc_0_sequencer_csr_writedata;    // mm_interconnect_1:modular_adc_0_sequencer_csr_writedata -> modular_adc_0:sequencer_csr_writedata
	wire   [0:0] mm_interconnect_1_modular_adc_0_sequencer_csr_address;      // mm_interconnect_1:modular_adc_0_sequencer_csr_address -> modular_adc_0:sequencer_csr_address
	wire         mm_interconnect_1_modular_adc_0_sequencer_csr_write;        // mm_interconnect_1:modular_adc_0_sequencer_csr_write -> modular_adc_0:sequencer_csr_write
	wire         mm_interconnect_1_modular_adc_0_sequencer_csr_read;         // mm_interconnect_1:modular_adc_0_sequencer_csr_read -> modular_adc_0:sequencer_csr_read
	wire  [31:0] mm_interconnect_1_modular_adc_0_sequencer_csr_readdata;     // modular_adc_0:sequencer_csr_readdata -> mm_interconnect_1:modular_adc_0_sequencer_csr_readdata
	wire  [31:0] mm_interconnect_1_modular_adc_0_sample_store_csr_writedata; // mm_interconnect_1:modular_adc_0_sample_store_csr_writedata -> modular_adc_0:sample_store_csr_writedata
	wire   [6:0] mm_interconnect_1_modular_adc_0_sample_store_csr_address;   // mm_interconnect_1:modular_adc_0_sample_store_csr_address -> modular_adc_0:sample_store_csr_address
	wire         mm_interconnect_1_modular_adc_0_sample_store_csr_write;     // mm_interconnect_1:modular_adc_0_sample_store_csr_write -> modular_adc_0:sample_store_csr_write
	wire         mm_interconnect_1_modular_adc_0_sample_store_csr_read;      // mm_interconnect_1:modular_adc_0_sample_store_csr_read -> modular_adc_0:sample_store_csr_read
	wire  [31:0] mm_interconnect_1_modular_adc_0_sample_store_csr_readdata;  // modular_adc_0:sample_store_csr_readdata -> mm_interconnect_1:modular_adc_0_sample_store_csr_readdata
	wire  [31:0] nios2_gen2_0_irq_irq;                                       // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         irq_mapper_receiver0_irq;                                   // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                              // systimer:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                   // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                          // jtag_uart:av_irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                   // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                          // modular_adc_0:sample_store_irq_irq -> irq_synchronizer_002:receiver_irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:onchip_flash_0_nreset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_flash_0:reset_n, rst_translator:in_reset, sdram:reset_n]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                     // nios2_gen2_0:jtag_debug_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [mm_interconnect_0:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, onchip_memory2_0:reset]
	wire         rst_controller_001_reset_out_reset_req;                     // rst_controller_001:reset_req -> onchip_memory2_0:reset_req
	wire         rst_controller_002_reset_out_reset;                         // rst_controller_002:reset_out -> [gpio:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, jtag_uart:rst_n, led:reset_n, mm_interconnect_0:peripheral_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_1:peripheral_bridge_reset_reset_bridge_in_reset_reset, modular_adc_0:reset_sink_reset_n, peripheral_bridge:reset, sysid:reset_n, systimer:reset_n]

	testcore_nios2_gen2_0 nios2_gen2_0 (
		.clk                                  (clk100_clk),                                                 //                       clk.clk
		.reset_n                              (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                            (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                            (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                         (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                               (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                           (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                        (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                              (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                          (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                      (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.jtag_debug_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                            (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                               (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                           (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                        (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                      (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                  (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.jtag_debug_resetrequest              (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.jtag_debug_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.jtag_debug_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.jtag_debug_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.jtag_debug_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.jtag_debug_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.jtag_debug_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.jtag_debug_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.jtag_debug_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                        ()                                                            // custom_instruction_master.readra
	);

	testcore_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk100_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)            //       .reset_req
	);

	altera_onchip_flash #(
		.INIT_FILENAME               (""),
		.INIT_FILENAME_SIM           (""),
		.DEVICE_FAMILY               ("MAX 10 FPGA"),
		.PART_NAME                   ("10M08SAE144C8GES"),
		.DEVICE_ID                   ("08"),
		.SECTOR1_START_ADDR          (512),
		.SECTOR1_END_ADDR            (4607),
		.SECTOR2_START_ADDR          (4608),
		.SECTOR2_END_ADDR            (8703),
		.SECTOR3_START_ADDR          (0),
		.SECTOR3_END_ADDR            (0),
		.SECTOR4_START_ADDR          (0),
		.SECTOR4_END_ADDR            (0),
		.SECTOR5_START_ADDR          (0),
		.SECTOR5_END_ADDR            (0),
		.MIN_VALID_ADDR              (512),
		.MAX_VALID_ADDR              (8703),
		.MIN_UFM_VALID_ADDR          (512),
		.MAX_UFM_VALID_ADDR          (8703),
		.AVMM_DATA_ADDR_WIDTH        (13),
		.AVMM_DATA_BURSTCOUNT_WIDTH  (4),
		.SECTOR_READ_PROTECTION_MODE (28),
		.FLASH_SEQ_READ_DATA_COUNT   (2),
		.FLASH_ADDR_ALIGNMENT_BITS   (1),
		.FLASH_READ_CYCLE_MAX_INDEX  (3),
		.FLASH_RESET_CYCLE_MAX_INDEX (25),
		.READ_AND_WRITE_MODE         (1),
		.WRAPPING_BURST_MODE         (0),
		.IS_DUAL_BOOT                ("False")
	) onchip_flash_0 (
		.clock                   (clk100_clk),                                          //    clk.clk
		.reset_n                 (~rst_controller_reset_out_reset),                     // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_onchip_flash_0_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_onchip_flash_0_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_0_onchip_flash_0_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_0_onchip_flash_0_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_0_onchip_flash_0_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_onchip_flash_0_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_onchip_flash_0_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_onchip_flash_0_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_1_onchip_flash_0_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_1_onchip_flash_0_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_1_onchip_flash_0_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_1_onchip_flash_0_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_1_onchip_flash_0_csr_readdata)        //       .readdata
	);

	testcore_sysid sysid (
		.clock    (clk40_clk),                                      //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	testcore_systimer systimer (
		.clk        (clk40_clk),                                //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.address    (mm_interconnect_1_systimer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_systimer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_systimer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_systimer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_systimer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)             //   irq.irq
	);

	testcore_jtag_uart jtag_uart (
		.clk            (clk40_clk),                                                 //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_001_receiver_irq)                          //               irq.irq
	);

	testcore_led led (
		.clk        (clk40_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	testcore_gpio gpio (
		.clk        (clk40_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_1_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_gpio_s1_readdata),   //                    .readdata
		.bidir_port (gpio_export)                           // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (16),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) peripheral_bridge (
		.clk              (clk40_clk),                                            //   clk.clk
		.reset            (rst_controller_002_reset_out_reset),                   // reset.reset
		.s0_waitrequest   (mm_interconnect_0_peripheral_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_peripheral_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_peripheral_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_peripheral_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_peripheral_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_peripheral_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_peripheral_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_peripheral_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_peripheral_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_peripheral_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (peripheral_bridge_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (peripheral_bridge_m0_readdata),                        //      .readdata
		.m0_readdatavalid (peripheral_bridge_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (peripheral_bridge_m0_burstcount),                      //      .burstcount
		.m0_writedata     (peripheral_bridge_m0_writedata),                       //      .writedata
		.m0_address       (peripheral_bridge_m0_address),                         //      .address
		.m0_write         (peripheral_bridge_m0_write),                           //      .write
		.m0_read          (peripheral_bridge_m0_read),                            //      .read
		.m0_byteenable    (peripheral_bridge_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (peripheral_bridge_m0_debugaccess)                      //      .debugaccess
	);

	testcore_sdram sdram (
		.clk            (clk100_clk),                               //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdr_addr),                                 //  wire.export
		.zs_ba          (sdr_ba),                                   //      .export
		.zs_cas_n       (sdr_cas_n),                                //      .export
		.zs_cke         (sdr_cke),                                  //      .export
		.zs_cs_n        (sdr_cs_n),                                 //      .export
		.zs_dq          (sdr_dq),                                   //      .export
		.zs_dqm         (sdr_dqm),                                  //      .export
		.zs_ras_n       (sdr_ras_n),                                //      .export
		.zs_we_n        (sdr_we_n)                                  //      .export
	);

	testcore_modular_adc_0 modular_adc_0 (
		.clock_clk                  (clk40_clk),                                                  //            clock.clk
		.reset_sink_reset_n         (~rst_controller_002_reset_out_reset),                        //       reset_sink.reset_n
		.adc_pll_clock_clk          (clk40_clk),                                                  //    adc_pll_clock.clk
		.adc_pll_locked_export      (adc_pll_locked_export),                                      //   adc_pll_locked.export
		.sequencer_csr_address      (mm_interconnect_1_modular_adc_0_sequencer_csr_address),      //    sequencer_csr.address
		.sequencer_csr_read         (mm_interconnect_1_modular_adc_0_sequencer_csr_read),         //                 .read
		.sequencer_csr_write        (mm_interconnect_1_modular_adc_0_sequencer_csr_write),        //                 .write
		.sequencer_csr_writedata    (mm_interconnect_1_modular_adc_0_sequencer_csr_writedata),    //                 .writedata
		.sequencer_csr_readdata     (mm_interconnect_1_modular_adc_0_sequencer_csr_readdata),     //                 .readdata
		.sample_store_csr_address   (mm_interconnect_1_modular_adc_0_sample_store_csr_address),   // sample_store_csr.address
		.sample_store_csr_read      (mm_interconnect_1_modular_adc_0_sample_store_csr_read),      //                 .read
		.sample_store_csr_write     (mm_interconnect_1_modular_adc_0_sample_store_csr_write),     //                 .write
		.sample_store_csr_writedata (mm_interconnect_1_modular_adc_0_sample_store_csr_writedata), //                 .writedata
		.sample_store_csr_readdata  (mm_interconnect_1_modular_adc_0_sample_store_csr_readdata),  //                 .readdata
		.sample_store_irq_irq       (irq_synchronizer_002_receiver_irq)                           // sample_store_irq.irq
	);

	testcore_mm_interconnect_0 mm_interconnect_0 (
		.clk_core_clk_clk                                    (clk100_clk),                                                 //                                  clk_core_clk.clk
		.clk_peri_clk_clk                                    (clk40_clk),                                                  //                                  clk_peri_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                             //      nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.onchip_memory2_0_reset1_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                         // onchip_memory2_0_reset1_reset_bridge_in_reset.reset
		.peripheral_bridge_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                         // peripheral_bridge_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                    (nios2_gen2_0_data_master_address),                           //                      nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                (nios2_gen2_0_data_master_waitrequest),                       //                                              .waitrequest
		.nios2_gen2_0_data_master_byteenable                 (nios2_gen2_0_data_master_byteenable),                        //                                              .byteenable
		.nios2_gen2_0_data_master_read                       (nios2_gen2_0_data_master_read),                              //                                              .read
		.nios2_gen2_0_data_master_readdata                   (nios2_gen2_0_data_master_readdata),                          //                                              .readdata
		.nios2_gen2_0_data_master_readdatavalid              (nios2_gen2_0_data_master_readdatavalid),                     //                                              .readdatavalid
		.nios2_gen2_0_data_master_write                      (nios2_gen2_0_data_master_write),                             //                                              .write
		.nios2_gen2_0_data_master_writedata                  (nios2_gen2_0_data_master_writedata),                         //                                              .writedata
		.nios2_gen2_0_data_master_debugaccess                (nios2_gen2_0_data_master_debugaccess),                       //                                              .debugaccess
		.nios2_gen2_0_instruction_master_address             (nios2_gen2_0_instruction_master_address),                    //               nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest         (nios2_gen2_0_instruction_master_waitrequest),                //                                              .waitrequest
		.nios2_gen2_0_instruction_master_read                (nios2_gen2_0_instruction_master_read),                       //                                              .read
		.nios2_gen2_0_instruction_master_readdata            (nios2_gen2_0_instruction_master_readdata),                   //                                              .readdata
		.nios2_gen2_0_instruction_master_readdatavalid       (nios2_gen2_0_instruction_master_readdatavalid),              //                                              .readdatavalid
		.nios2_gen2_0_debug_mem_slave_address                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //                  nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                  (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                              .write
		.nios2_gen2_0_debug_mem_slave_read                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                              .read
		.nios2_gen2_0_debug_mem_slave_readdata               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                              .readdata
		.nios2_gen2_0_debug_mem_slave_writedata              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                              .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                              .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                              .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                              .debugaccess
		.onchip_flash_0_data_address                         (mm_interconnect_0_onchip_flash_0_data_address),              //                           onchip_flash_0_data.address
		.onchip_flash_0_data_write                           (mm_interconnect_0_onchip_flash_0_data_write),                //                                              .write
		.onchip_flash_0_data_read                            (mm_interconnect_0_onchip_flash_0_data_read),                 //                                              .read
		.onchip_flash_0_data_readdata                        (mm_interconnect_0_onchip_flash_0_data_readdata),             //                                              .readdata
		.onchip_flash_0_data_writedata                       (mm_interconnect_0_onchip_flash_0_data_writedata),            //                                              .writedata
		.onchip_flash_0_data_burstcount                      (mm_interconnect_0_onchip_flash_0_data_burstcount),           //                                              .burstcount
		.onchip_flash_0_data_readdatavalid                   (mm_interconnect_0_onchip_flash_0_data_readdatavalid),        //                                              .readdatavalid
		.onchip_flash_0_data_waitrequest                     (mm_interconnect_0_onchip_flash_0_data_waitrequest),          //                                              .waitrequest
		.onchip_memory2_0_s1_address                         (mm_interconnect_0_onchip_memory2_0_s1_address),              //                           onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                           (mm_interconnect_0_onchip_memory2_0_s1_write),                //                                              .write
		.onchip_memory2_0_s1_readdata                        (mm_interconnect_0_onchip_memory2_0_s1_readdata),             //                                              .readdata
		.onchip_memory2_0_s1_writedata                       (mm_interconnect_0_onchip_memory2_0_s1_writedata),            //                                              .writedata
		.onchip_memory2_0_s1_byteenable                      (mm_interconnect_0_onchip_memory2_0_s1_byteenable),           //                                              .byteenable
		.onchip_memory2_0_s1_chipselect                      (mm_interconnect_0_onchip_memory2_0_s1_chipselect),           //                                              .chipselect
		.onchip_memory2_0_s1_clken                           (mm_interconnect_0_onchip_memory2_0_s1_clken),                //                                              .clken
		.peripheral_bridge_s0_address                        (mm_interconnect_0_peripheral_bridge_s0_address),             //                          peripheral_bridge_s0.address
		.peripheral_bridge_s0_write                          (mm_interconnect_0_peripheral_bridge_s0_write),               //                                              .write
		.peripheral_bridge_s0_read                           (mm_interconnect_0_peripheral_bridge_s0_read),                //                                              .read
		.peripheral_bridge_s0_readdata                       (mm_interconnect_0_peripheral_bridge_s0_readdata),            //                                              .readdata
		.peripheral_bridge_s0_writedata                      (mm_interconnect_0_peripheral_bridge_s0_writedata),           //                                              .writedata
		.peripheral_bridge_s0_burstcount                     (mm_interconnect_0_peripheral_bridge_s0_burstcount),          //                                              .burstcount
		.peripheral_bridge_s0_byteenable                     (mm_interconnect_0_peripheral_bridge_s0_byteenable),          //                                              .byteenable
		.peripheral_bridge_s0_readdatavalid                  (mm_interconnect_0_peripheral_bridge_s0_readdatavalid),       //                                              .readdatavalid
		.peripheral_bridge_s0_waitrequest                    (mm_interconnect_0_peripheral_bridge_s0_waitrequest),         //                                              .waitrequest
		.peripheral_bridge_s0_debugaccess                    (mm_interconnect_0_peripheral_bridge_s0_debugaccess),         //                                              .debugaccess
		.sdram_s1_address                                    (mm_interconnect_0_sdram_s1_address),                         //                                      sdram_s1.address
		.sdram_s1_write                                      (mm_interconnect_0_sdram_s1_write),                           //                                              .write
		.sdram_s1_read                                       (mm_interconnect_0_sdram_s1_read),                            //                                              .read
		.sdram_s1_readdata                                   (mm_interconnect_0_sdram_s1_readdata),                        //                                              .readdata
		.sdram_s1_writedata                                  (mm_interconnect_0_sdram_s1_writedata),                       //                                              .writedata
		.sdram_s1_byteenable                                 (mm_interconnect_0_sdram_s1_byteenable),                      //                                              .byteenable
		.sdram_s1_readdatavalid                              (mm_interconnect_0_sdram_s1_readdatavalid),                   //                                              .readdatavalid
		.sdram_s1_waitrequest                                (mm_interconnect_0_sdram_s1_waitrequest),                     //                                              .waitrequest
		.sdram_s1_chipselect                                 (mm_interconnect_0_sdram_s1_chipselect)                       //                                              .chipselect
	);

	testcore_mm_interconnect_1 mm_interconnect_1 (
		.clk_core_clk_clk                                    (clk100_clk),                                                 //                                  clk_core_clk.clk
		.clk_peri_clk_clk                                    (clk40_clk),                                                  //                                  clk_peri_clk.clk
		.onchip_flash_0_nreset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                             //   onchip_flash_0_nreset_reset_bridge_in_reset.reset
		.peripheral_bridge_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                         // peripheral_bridge_reset_reset_bridge_in_reset.reset
		.peripheral_bridge_m0_address                        (peripheral_bridge_m0_address),                               //                          peripheral_bridge_m0.address
		.peripheral_bridge_m0_waitrequest                    (peripheral_bridge_m0_waitrequest),                           //                                              .waitrequest
		.peripheral_bridge_m0_burstcount                     (peripheral_bridge_m0_burstcount),                            //                                              .burstcount
		.peripheral_bridge_m0_byteenable                     (peripheral_bridge_m0_byteenable),                            //                                              .byteenable
		.peripheral_bridge_m0_read                           (peripheral_bridge_m0_read),                                  //                                              .read
		.peripheral_bridge_m0_readdata                       (peripheral_bridge_m0_readdata),                              //                                              .readdata
		.peripheral_bridge_m0_readdatavalid                  (peripheral_bridge_m0_readdatavalid),                         //                                              .readdatavalid
		.peripheral_bridge_m0_write                          (peripheral_bridge_m0_write),                                 //                                              .write
		.peripheral_bridge_m0_writedata                      (peripheral_bridge_m0_writedata),                             //                                              .writedata
		.peripheral_bridge_m0_debugaccess                    (peripheral_bridge_m0_debugaccess),                           //                                              .debugaccess
		.gpio_s1_address                                     (mm_interconnect_1_gpio_s1_address),                          //                                       gpio_s1.address
		.gpio_s1_write                                       (mm_interconnect_1_gpio_s1_write),                            //                                              .write
		.gpio_s1_readdata                                    (mm_interconnect_1_gpio_s1_readdata),                         //                                              .readdata
		.gpio_s1_writedata                                   (mm_interconnect_1_gpio_s1_writedata),                        //                                              .writedata
		.gpio_s1_chipselect                                  (mm_interconnect_1_gpio_s1_chipselect),                       //                                              .chipselect
		.jtag_uart_avalon_jtag_slave_address                 (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),      //                   jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),        //                                              .write
		.jtag_uart_avalon_jtag_slave_read                    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),         //                                              .read
		.jtag_uart_avalon_jtag_slave_readdata                (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),     //                                              .readdata
		.jtag_uart_avalon_jtag_slave_writedata               (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),    //                                              .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest             (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest),  //                                              .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect              (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),   //                                              .chipselect
		.led_s1_address                                      (mm_interconnect_1_led_s1_address),                           //                                        led_s1.address
		.led_s1_write                                        (mm_interconnect_1_led_s1_write),                             //                                              .write
		.led_s1_readdata                                     (mm_interconnect_1_led_s1_readdata),                          //                                              .readdata
		.led_s1_writedata                                    (mm_interconnect_1_led_s1_writedata),                         //                                              .writedata
		.led_s1_chipselect                                   (mm_interconnect_1_led_s1_chipselect),                        //                                              .chipselect
		.modular_adc_0_sample_store_csr_address              (mm_interconnect_1_modular_adc_0_sample_store_csr_address),   //                modular_adc_0_sample_store_csr.address
		.modular_adc_0_sample_store_csr_write                (mm_interconnect_1_modular_adc_0_sample_store_csr_write),     //                                              .write
		.modular_adc_0_sample_store_csr_read                 (mm_interconnect_1_modular_adc_0_sample_store_csr_read),      //                                              .read
		.modular_adc_0_sample_store_csr_readdata             (mm_interconnect_1_modular_adc_0_sample_store_csr_readdata),  //                                              .readdata
		.modular_adc_0_sample_store_csr_writedata            (mm_interconnect_1_modular_adc_0_sample_store_csr_writedata), //                                              .writedata
		.modular_adc_0_sequencer_csr_address                 (mm_interconnect_1_modular_adc_0_sequencer_csr_address),      //                   modular_adc_0_sequencer_csr.address
		.modular_adc_0_sequencer_csr_write                   (mm_interconnect_1_modular_adc_0_sequencer_csr_write),        //                                              .write
		.modular_adc_0_sequencer_csr_read                    (mm_interconnect_1_modular_adc_0_sequencer_csr_read),         //                                              .read
		.modular_adc_0_sequencer_csr_readdata                (mm_interconnect_1_modular_adc_0_sequencer_csr_readdata),     //                                              .readdata
		.modular_adc_0_sequencer_csr_writedata               (mm_interconnect_1_modular_adc_0_sequencer_csr_writedata),    //                                              .writedata
		.onchip_flash_0_csr_address                          (mm_interconnect_1_onchip_flash_0_csr_address),               //                            onchip_flash_0_csr.address
		.onchip_flash_0_csr_write                            (mm_interconnect_1_onchip_flash_0_csr_write),                 //                                              .write
		.onchip_flash_0_csr_read                             (mm_interconnect_1_onchip_flash_0_csr_read),                  //                                              .read
		.onchip_flash_0_csr_readdata                         (mm_interconnect_1_onchip_flash_0_csr_readdata),              //                                              .readdata
		.onchip_flash_0_csr_writedata                        (mm_interconnect_1_onchip_flash_0_csr_writedata),             //                                              .writedata
		.sysid_control_slave_address                         (mm_interconnect_1_sysid_control_slave_address),              //                           sysid_control_slave.address
		.sysid_control_slave_readdata                        (mm_interconnect_1_sysid_control_slave_readdata),             //                                              .readdata
		.systimer_s1_address                                 (mm_interconnect_1_systimer_s1_address),                      //                                   systimer_s1.address
		.systimer_s1_write                                   (mm_interconnect_1_systimer_s1_write),                        //                                              .write
		.systimer_s1_readdata                                (mm_interconnect_1_systimer_s1_readdata),                     //                                              .readdata
		.systimer_s1_writedata                               (mm_interconnect_1_systimer_s1_writedata),                    //                                              .writedata
		.systimer_s1_chipselect                              (mm_interconnect_1_systimer_s1_chipselect)                    //                                              .chipselect
	);

	testcore_irq_mapper irq_mapper (
		.clk           (clk100_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk40_clk),                          //       receiver_clk.clk
		.sender_clk     (clk100_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk40_clk),                          //       receiver_clk.clk
		.sender_clk     (clk100_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk40_clk),                          //       receiver_clk.clk
		.sender_clk     (clk100_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk100_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk100_clk),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk40_clk),                          //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
